b0VIM 8.0      9 I]#   root                                    suram-VirtualBox                        ~root/youngeun/Server_Thread.java                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            utf-8U3210    #"! U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 tp	           r                     ��������|       s                            �                     \       �              ��������L       N             ��������J       �             ��������L       �             ��������o       0             ��������q       �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     ad          r       �  �  �  �  t  b  O  3     �  �  �  �  �  �  �  �  �  q  ]  L  *      �  �  �  �  �  �  �  �  �  �  �  \    �  �  �  |  X    �  �  �  �  v  u  e  L  A    �
  �
  b
  )
  
  �	  �	  U	  	  �  �  �  w  L    �  �  �  �  [  5    �  �  �  �  |  ]  ?      �  �  �  u  W  K  3    �  �  �  �  �  T  $    �  �  �  �  R  4    �  �  �  m  A                                        		                 break;		  				 System.out.println(result); 		                 oos.writeObject(result); 		                 result=selectDB_str(2,id); 		                 id=(String)ois.readObject(); 		                 String id=new String(); 		       case "temp_message_count": 		                 break; 				 oos.writeObject(result); 		                 System.out.println(result); 		                 result=selectDB_str(1,""); 		       case "lately_mid": 		                 break; 				 System.out.println(result); 				 oos.writeObject(result); 		                 result=selectDB_str(0,p_id); 		                 p_id=(String)ois.readObject(); 		                 String p_id=new String(); 		       case "get_mid": 				 break; 				 sendTK(0,token); 				 token=(String)ois.readObject(); 				 String token=new String(); 			case "update token": 				 break; 				 oos.writeObject(result); 				 result= selectDB(5,gData); 				 gData=(CommentRequest)ois.readObject(); 				 CommentRequest gData=new CommentRequest(); 			case "get_info": 				 break; 				 System.out.println("datalist:"+result); 				 oos.writeObject(result); 				 result=selectDB(4,lData); 				 lData=(loginData)ois.readObject(); 			         loginData lData=new loginData(); 			case "login": 				 break; 				 System.out.println(obj_result); 				 oos.writeObject(obj_result); 				 obj_result=selectDB_obj(0,s_id); 				 System.out.println("get_messge's s_id:"+s_id); 				 s_id=(String)ois.readObject(); 				 String s_id=new String(); 		        case "get_message":                                  break;                                  insertDB(2,mData); 				 mData=(messageData)ois.readObject();	 				 messageData mData=new messageData(); 			case "send_message":                                  break;                                 oos.writeObject(result);                                 result=selectDB(1,rData2); 			       rData2=(CommentRequest)ois.readObject();                                CommentRequest rData2=new CommentRequest();                         case "choose_comment":                                 break;                                 oos.writeObject(result);                                 result=selectDB(0,rData);                                 rData=(CommentRequest)ois.readObject(); 				CommentRequest rData=new CommentRequest();                         case "today_comment": 				break; 				//messageTab setting 			case "init":                  switch(type){                 String input="";                 ArrayList<String> inputs=new ArrayList<>();              System.out.println(type);            // ArrayList<String> result=new ArrayList<String>(); 	    type=(String)ois.readObject(); 	    try{              ObjectOutputStream oos = new ObjectOutputStream(outputStream);             OutputStream outputStream = client.getOutputStream();             ObjectInputStream ois = new ObjectInputStream(inputStream);             InputStream inputStream = client.getInputStream();             System.out.println("make client!");    	    try{              public void run(){      }      	type="";         this.client=socket;     Server_Thread(Socket socket){ 	int int_result; 	String str_result; 	ArrayList<Object> obj_result; 	ArrayList<String> result; 	String type = ""; 	Socket client;  public class Server_Thread extends Thread{    import java.text.SimpleDateFormat; import java.sql.*; import java.util.ArrayList; import java.net.*; import java.io.*; import com.example.youngeun.parentapp.*; import java.util.Date; import java.text.SimpleDateFormat;  package com.example.youngeun.parentapp; ad  O  /     q       �  �  [      �  �  �  �  Z  &  �  p    �  �  �  l  B  A  /    �  �  �  �  �  l  f  >    �
  �
  i
  \
  9
  2
  &
  
  
   
  �	  �	  �	  �	  �	  �	  	  W	  >	  '	  	  �  �  �  �  �  �  ^  �  �  �  �  �  �  �  �  �  @  !         �  �  �  w  p  j  i  �  �  �  �  B  �  �  �  Y  *  "    �  �  �  �  �  �  �  �  �  ~  y  x  a  I  F  A  ;  7  6  1  /  .                                                                                                                                                                                                                                                                                                                                                 }               }      		 		e.printStackTrace();} 		}catch(Exception e){  			} 			    			                                   break; 			                                    pstmt.executeUpdate();   				  } 				     pstmt.setInt(6,0); 				  else{ 				  } 		                     pstmt.setInt(6,1);			   				  if((mData.getState()).equals("final")){	 				  pstmt.setString(5,mData.getRequest());                                   pstmt.setString(4,mData.getP_id());                                   pstmt.setString(3,mData.getMdate());                                   pstmt.setString(2,mData.getMessage()); 				  pstmt.setString(1,mData.getM_id()); 				  pstmt=conn.prepareStatement(sql); 				  		        	  sql="insert into message_tbl(m_id,m_cont,m_date,p_id,m_req,final) values(?,?,?,?,?,?);";                                  				} 					} 						stmt.executeUpdate(sql); 						sql="delete from message_tbl where m_id='"+mData.getM_id()+"';"; 					 					if((rs.getInt("count(*)"))!=0){ 				 				if(rs.next()){  				rs=stmt.executeQuery(sql); 				sql="select count(*) from message_tbl where m_id='"+mData.getM_id()+"';";  				messageData mData= (messageData)object; 				case 2: 			 			switch(type){   			stmt=conn.createStatement(); 					"jdbc:mysql://localhost/tidsnotedb?characterEncoding=UTF-8"+"&user=suram&password=suram"); 			conn=DriverManager.getConnection( 			Class.forName("com.mysql.cj.jdbc.Driver");  		try { 	 		ArrayList<String> datalist=new ArrayList<String>(); 		String sql = ""; 		PreparedStatement pstmt = null; 		ResultSet rs = null; 		Statement stmt = null;                 Connection conn = null;          public static void insertDB(int type,Object object ){     }      		  return datalist;  			       	e.printStackTrace();} 			}catch(Exception e){  			}//switch 					break; 					} 					       datalist.add(tempMSG); 					        					       tempMSG.setM_id(rs.getString("m_id")); 					       tempMSG.setRequest(rs.getString("m_req")); 					       tempMSG.setMessage(rs.getString("m_cont")); 					       tempMSG.setP_id(rs.getString("p_id")); 					       tempMSG=new messageData();	 					 					if(rs.next()){  					messageData tempMSG;  					rs=stmt.executeQuery(sql); 					sql="select * from message_tbl where final=0 and p_id='"+p_id2+"';"; 				        String p_id2=(String)string; 			       case 1:                                     break;                                     }//while                                             datalist.add(messagedata);  					    messagedata.setM_id(rs.getString("m_id"));                                             messagedata.setRequest(rs.getString("m_req"));                                             messagedata.setMessage(rs.getString("m_cont"));                                             messagedata.setMdate(rs.getString("m_date")); 					    messagedata.setP_id(rs.getString("p_id"));                                             messagedata= new messageData();                                      while(rs.next()){                                      messageData messagedata;                                      rs=stmt.executeQuery(sql);                                     sql="select * from message_tbl where final=1 and p_id='"+s_id+"' order by m_id desc"; 					  } 						s_id=rs2.getString("p_id"); ad  0  \            �  �  �  \  \  �  �  �  �  �  �  s  r  \  V        �  �  �  �  T  @  ?  5  /  �  |  Y  X  D  >  6     �  �  �  A    �
  �
  f
  e
  d
  
  �	  �	  �	  p	  	  �  �  �  �  N      �  �  ~  H    �  �  L  B    �  �  V  U  !  �  �  i  h  �  �  �  �  /  �  �  �  �  �  �  �  ~  z  W  $  �  �  �      				   // String t_name=rs.getString("t_name"); 				    String date=rs.getString("c_date"); 				    String name=rs.getString("s_name"); 			           // String s_id=rs.getString("s_id"); 				 if (rs.getInt("final")!=0){	  			 				 }else{ //교사가 코멘트를 작성했을 경우  					   break;                                     }                                             datalist.add(t_name);                                             String t_name=rs3.getString("c_name");                                     if(rs3.next()){                                    rs3=stmt.executeQuery(sql);                                  sql="select c_name from class_tbl,comment_tbl where s_id='"+rData.getS_id()+"';";                                   }                                             datalist.add(t_name);                                             String t_name=rs2.getString("t_name");                                     if(rs2.next()){                                      rs2=stmt.executeQuery(sql);                                      sql=sql+"(select t_id from student_tbl where s_id='"+rData.getS_id()+"');"; 				     sql="select t_name from teacher_tbl where t_id="; 				   }                                      datalist.add("");                                     datalist.add(" 작성되지 않았습니다.");                                    // datalist.add(m_menu);                                     datalist.add("");                                     datalist.add("");                                     datalist.add(""); 				        datalist.add(date);                                         datalist.add(name); 					    					   String date=simpleformat.format(new Date()); 					   SimpleDateFormat simpleformat=new SimpleDateFormat("yyyy-MM-dd"); 					   String name=rs4.getString("s_name"); 				   if(rs4.next()){                                      rs4=stmt.executeQuery(sql);                                     sql=sql+"where S.s_id='"+rData.getS_id()+"';";                                     sql=sql+" from student_tbl S "; 					    sql="select S.s_name"; 				     					   System.out.println("today's comment not yet.."); 				    if(!rs.next()){//교사가 코멘트를 작성하지 않았을 경우   				    rs=stmt.executeQuery(sql); 				    sql=sql+" C.c_date>CURRENT_DATE();";//m_menu  				    sql=sql+"where C.s_id='"+rData.getS_id()+"' and S.s_id=C.s_id and"; 				    sql=sql+" from student_tbl S,comment_tbl C "; 		                    sql=sql+"C.c_feel,C.c_meal,C.c_health,C.c_comment,C.c_same"; 				    sql="select C.final,S.s_name,C.c_date,"; 	     				    CommentRequest rData=(CommentRequest)object; 			    case 0://코멘트 조회(새로고침)-당일 			     		    		    switch(type){  		    stmt=conn.createStatement(); 		    conn=DriverManager.getConnection("jdbc:mysql://localhost/tidsnotedb?characterEncoding=UTF-8"+"&user=suram&password=suram"); 		    Class.forName("com.mysql.cj.jdbc.Driver"); 	     	    try{  	    String sql=""; 	    ArrayList<String> datalist=new ArrayList<>(); 	    PreparedStatement pstmt=null; 	    ResultSet rs,rs2,rs3,rs4,rs5=null; 	    Statement stmt=null; 	    Connection conn=null;             public static ArrayList<String> selectDB(int type, Object object){     } 	    return datalist;              }                     e.printStackTrace(); 	    }catch(Exception e){ 		    }                                      break;		                                         }                                          datalist.add(rs					    String str_count=rs.getInt("count(*)");                                     if(rs.next()){                                      rs=stmt.executeQuery(sql); ad  �   '     \       �  �  X  W  O  5    �  �  �  �  �  �  �  w  ]  5    �  �  �  �  �  �    �  �  �  �  �  �  V  P    �  �  J    �
  �
  �
  �
  h
  _
  ?
  �	  �	  h	  g	  P	  #	  �  �  �  _  ?  	  �  �  a    �  �  �  "  !  �  �  �  Y    �  �  �  B  A    �  x  U  T  S  R  C  B  	    �  �  �  W  '                                                                                                                                                                 				   // String t_name=rs.getString("t_name"); 				    String date=rs.getString("c_date"); 				    String name=rs.getString("s_name"); 			           // String s_id=rs.getString("s_id"); 				 if (rs.getInt("final")!=0){	  			 				 }else{ //교사가 코멘트를 작성했을 경우  					   break;                                     }                                             datalist.add(t_name);                                             String t_name=rs3.getString("c_name");                                     if(rs3.next()){                                    rs3=stmt.executeQuery(sql);                                  sql="select c_name from class_tbl,comment_tbl where s_id='"+rData.getS_id()+"';";                                   }                                             datalist.add(t_name);                                             String t_name=rs2.getString("t_name");                                     if(rs2.next()){                                      rs2=stmt.executeQuery(sql);                                      sql=sql+"(select t_id from student_tbl where s_id='"+rData.getS_id()+"');"; 				     sql="select t_name from teacher_tbl where t_id="; 				   }                                      datalist.add("");                                     datalist.add(" 작성되지 않았습니다.");                                    // datalist.add(m_menu);                                     datalist.add("");                                     datalist.add("");                                     datalist.add(""); 				        datalist.add(date);                                         datalist.add(name); 					    					   String date=simpleformat.format(new Date()); 					   SimpleDateFormat simpleformat=new SimpleDateFormat("yyyy-MM-dd"); 					   String name=rs4.getString("s_name"); 				   if(rs4.next()){                                      rs4=stmt.executeQuery(sql);                                     sql=sql+"where S.s_id='"+rData.getS_id()+"';";                                     sql=sql+" from student_tbl S "; 					    sql="select S.s_name"; 				     					   System.out.println("today's comment not yet.."); 				    if(!rs.next()){//교사가 코멘트를 작성하지 않았을 경우   				    rs=stmt.executeQuery(sql); 				    sql=sql+" C.c_date>CURRENT_DATE();";//m_menu  				    sql=sql+"where C.s_id='"+rData.getS_id()+"' and S.s_id=C.s_id and"; 				    sql=sql+" from student_tbl S,comment_tbl C "; 		                    sql=sql+"C.c_feel,C.c_meal,C.c_health,C.c_comment,C.c_same"; 				    sql="select C.final,S.s_name,C.c_date,"; 	     				    CommentRequest rData=(CommentRequest)object; 			    case 0://코멘트 조회(새로고침)-당일 			     		    		    switch(type){  		    stmt=conn.createStatement(); 		    conn=DriverManager.getConnection("jdbc:mysql://localhost/tidsnotedb?characterEncoding=UTF-8"+"&user=suram&password=suram"); 		    Class.forName("com.mysql.cj.jdbc.Driver"); 	     	    try{  	    String sql=""; 	    ArrayList<String> datalist=new ArrayList<>(); 	    PreparedStatement pstmt=null; 	    ResultSet rs,rs2,rs3,rs4,rs5=null; 	    Statement stmt=null; 	    Connection conn=null;             public static ArrayList<String> selectDB(int type, Object object){     } 	    return datalist;              }                     e.printStackTrace(); 	    }catch(Exception e){ 		    }                                      break;		                                         }                                          datalist.add(rs.getString("count(*)")); 